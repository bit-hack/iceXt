/*     _          _  ________
 *    (_)_______ | |/ /_  __/
 *   / / ___/ _ \|   / / /
 *  / / /__/  __/   | / /
 * /_/\___/\___/_/|_|/_/
 *
**/

`ifdef INCLUDE_CONFIG_VH
`define INCLUDE_CONFIG_VH

//`define CFG_ADLIB_ENABLE

`endif
