`ifdef INCLUDE_CONFIG_VH
`define INCLUDE_CONFIG_VH

//`define CFG_ADLIB_ENABLE

`endif
